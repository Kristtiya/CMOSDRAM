magic
tech sky130A
timestamp 1614907382
<< nwell >>
rect -275 125 205 440
rect -20 10 205 125
<< nmos >>
rect -190 -65 -175 35
rect -125 -65 -110 35
rect -185 -220 -170 -120
rect -200 -350 -140 -250
rect 50 -185 65 -85
rect 115 -185 130 -85
rect 80 -350 140 -250
<< pmos >>
rect -200 320 -140 420
rect -10 320 50 420
rect -195 145 -180 245
rect -130 145 -115 245
rect 30 190 45 290
rect 55 30 70 130
rect 120 30 135 130
<< ndiff >>
rect -240 20 -190 35
rect -240 -50 -225 20
rect -205 -50 -190 20
rect -240 -65 -190 -50
rect -175 20 -125 35
rect -175 -50 -160 20
rect -140 -50 -125 20
rect -175 -65 -125 -50
rect -110 20 -60 35
rect -110 -50 -95 20
rect -75 -50 -60 20
rect -110 -65 -60 -50
rect -235 -135 -185 -120
rect -235 -205 -220 -135
rect -200 -205 -185 -135
rect -235 -220 -185 -205
rect -170 -135 -120 -120
rect -170 -205 -155 -135
rect -135 -205 -120 -135
rect -170 -220 -120 -205
rect -250 -265 -200 -250
rect -250 -335 -235 -265
rect -215 -335 -200 -265
rect -250 -350 -200 -335
rect -140 -265 -95 -250
rect -140 -335 -130 -265
rect -110 -335 -95 -265
rect -140 -350 -95 -335
rect 0 -100 50 -85
rect 0 -170 15 -100
rect 35 -170 50 -100
rect 0 -185 50 -170
rect 65 -100 115 -85
rect 65 -170 80 -100
rect 100 -170 115 -100
rect 65 -185 115 -170
rect 130 -100 180 -85
rect 130 -170 145 -100
rect 165 -170 180 -100
rect 130 -185 180 -170
rect 30 -265 80 -250
rect 30 -335 45 -265
rect 65 -335 80 -265
rect 30 -350 80 -335
rect 140 -265 190 -250
rect 140 -335 155 -265
rect 175 -335 190 -265
rect 140 -350 190 -335
<< pdiff >>
rect -255 405 -200 420
rect -255 335 -240 405
rect -215 335 -200 405
rect -255 320 -200 335
rect -140 405 -90 420
rect -140 335 -125 405
rect -105 335 -90 405
rect -140 320 -90 335
rect -60 405 -10 420
rect -60 335 -45 405
rect -25 335 -10 405
rect -60 320 -10 335
rect 50 405 100 420
rect 50 335 65 405
rect 85 335 100 405
rect 50 320 100 335
rect -245 230 -195 245
rect -245 160 -230 230
rect -210 160 -195 230
rect -245 145 -195 160
rect -180 230 -130 245
rect -180 160 -165 230
rect -145 160 -130 230
rect -180 145 -130 160
rect -115 230 -65 245
rect -115 160 -100 230
rect -80 160 -65 230
rect -115 145 -65 160
rect -20 275 30 290
rect -20 205 -5 275
rect 15 205 30 275
rect -20 190 30 205
rect 45 275 95 290
rect 45 205 60 275
rect 80 205 95 275
rect 45 190 95 205
rect 5 115 55 130
rect 5 45 20 115
rect 40 45 55 115
rect 5 30 55 45
rect 70 115 120 130
rect 70 45 85 115
rect 105 45 120 115
rect 70 30 120 45
rect 135 115 185 130
rect 135 45 150 115
rect 170 45 185 115
rect 135 30 185 45
<< ndiffc >>
rect -225 -50 -205 20
rect -160 -50 -140 20
rect -95 -50 -75 20
rect -220 -205 -200 -135
rect -155 -205 -135 -135
rect -235 -335 -215 -265
rect -130 -335 -110 -265
rect 15 -170 35 -100
rect 80 -170 100 -100
rect 145 -170 165 -100
rect 45 -335 65 -265
rect 155 -335 175 -265
<< pdiffc >>
rect -240 335 -215 405
rect -125 335 -105 405
rect -45 335 -25 405
rect 65 335 85 405
rect -230 160 -210 230
rect -165 160 -145 230
rect -100 160 -80 230
rect -5 205 15 275
rect 60 205 80 275
rect 20 45 40 115
rect 85 45 105 115
rect 150 45 170 115
<< psubdiff >>
rect -120 -135 -70 -120
rect -120 -205 -105 -135
rect -85 -205 -70 -135
rect -120 -220 -70 -205
<< nsubdiff >>
rect 95 275 145 290
rect 95 205 110 275
rect 130 205 145 275
rect 95 190 145 205
<< psubdiffcont >>
rect -105 -205 -85 -135
<< nsubdiffcont >>
rect 110 205 130 275
<< poly >>
rect -200 420 -140 435
rect -10 420 50 435
rect 155 400 195 410
rect 155 380 165 400
rect 185 380 195 400
rect 155 370 195 380
rect -200 305 -140 320
rect -10 305 50 320
rect -155 300 -140 305
rect -155 295 -35 300
rect -155 285 -30 295
rect 30 290 45 305
rect -50 280 -30 285
rect -195 245 -180 260
rect -130 245 -115 260
rect -45 180 -30 280
rect 30 180 45 190
rect -45 165 45 180
rect 180 175 195 370
rect -195 90 -180 145
rect -130 130 -115 145
rect -130 120 -90 130
rect -130 100 -120 120
rect -100 100 -90 120
rect -130 90 -90 100
rect -195 80 -155 90
rect -195 60 -185 80
rect -165 60 -155 80
rect -195 50 -155 60
rect -190 35 -175 50
rect -125 35 -110 90
rect -190 -80 -175 -65
rect -125 -80 -110 -65
rect -45 -75 -30 165
rect 120 160 195 175
rect 55 130 70 145
rect 120 130 135 160
rect 55 -30 70 30
rect 120 10 135 30
rect 95 0 135 10
rect 95 -20 105 0
rect 125 -20 135 0
rect 95 -30 135 -20
rect 30 -40 70 -30
rect 30 -60 40 -40
rect 60 -60 70 -40
rect 30 -70 70 -60
rect -65 -90 -30 -75
rect 50 -85 65 -70
rect 115 -85 130 -30
rect -185 -120 -170 -105
rect -185 -235 -170 -220
rect -200 -250 -140 -235
rect -200 -365 -140 -350
rect -180 -390 -165 -365
rect -65 -390 -50 -90
rect 50 -200 65 -185
rect 115 -200 130 -185
rect -15 -210 25 -200
rect -15 -230 -5 -210
rect 15 -230 25 -210
rect -15 -240 25 -230
rect -10 -305 5 -240
rect 80 -250 140 -235
rect -25 -315 15 -305
rect -25 -335 -15 -315
rect 5 -335 15 -315
rect -25 -345 15 -335
rect 80 -365 140 -350
rect 80 -390 95 -365
rect -180 -400 -140 -390
rect -180 -420 -170 -400
rect -150 -420 -140 -400
rect -180 -430 -140 -420
rect -80 -400 -40 -390
rect -80 -420 -70 -400
rect -50 -420 -40 -400
rect -80 -430 -40 -420
rect 75 -400 115 -390
rect 75 -420 85 -400
rect 105 -420 115 -400
rect 75 -430 115 -420
<< polycont >>
rect 165 380 185 400
rect -120 100 -100 120
rect -185 60 -165 80
rect 105 -20 125 0
rect 40 -60 60 -40
rect -5 -230 15 -210
rect -15 -335 5 -315
rect -170 -420 -150 -400
rect -70 -420 -50 -400
rect 85 -420 105 -400
<< locali >>
rect -275 445 75 465
rect 55 415 75 445
rect 115 445 205 465
rect -250 410 -205 415
rect -275 405 -205 410
rect -275 390 -240 405
rect -250 335 -240 390
rect -215 335 -205 405
rect -250 325 -205 335
rect -135 405 -95 415
rect -135 335 -125 405
rect -105 335 -95 405
rect -135 325 -95 335
rect -55 405 -15 415
rect -55 335 -45 405
rect -25 335 -15 405
rect -55 325 -15 335
rect 55 405 95 415
rect 55 335 65 405
rect 85 335 95 405
rect 55 325 95 335
rect 115 330 135 445
rect 155 400 205 410
rect 155 380 165 400
rect 185 390 205 400
rect 185 380 195 390
rect 155 370 195 380
rect -135 280 -115 325
rect -55 300 -35 325
rect 115 310 180 330
rect -220 260 -115 280
rect -90 280 -35 300
rect -220 240 -200 260
rect -90 240 -70 280
rect -240 230 -200 240
rect -240 160 -230 230
rect -210 160 -200 230
rect -240 150 -200 160
rect -175 230 -135 240
rect -175 160 -165 230
rect -145 160 -135 230
rect -175 150 -135 160
rect -110 230 -70 240
rect -110 160 -100 230
rect -80 170 -70 230
rect -15 275 25 285
rect -15 205 -5 275
rect 15 205 25 275
rect -15 195 25 205
rect 50 275 140 285
rect 50 205 60 275
rect 80 205 110 275
rect 130 205 140 275
rect 50 195 140 205
rect 5 175 25 195
rect -80 160 -50 170
rect -110 150 -50 160
rect 5 155 110 175
rect -235 130 -215 150
rect -235 120 -90 130
rect -235 110 -120 120
rect -235 30 -215 110
rect -130 100 -120 110
rect -100 100 -90 120
rect -130 90 -90 100
rect -195 80 -155 90
rect -195 60 -185 80
rect -165 70 -155 80
rect -70 70 -50 150
rect 90 125 110 155
rect 160 125 180 310
rect -165 60 -50 70
rect -195 50 -50 60
rect 10 115 50 125
rect -90 30 -70 50
rect 10 45 20 115
rect 40 45 50 115
rect 10 35 50 45
rect 75 115 115 125
rect 75 45 85 115
rect 105 45 115 115
rect 75 35 115 45
rect 140 115 180 125
rect 140 45 150 115
rect 170 45 180 115
rect 140 35 180 45
rect -235 20 -195 30
rect -235 -40 -225 20
rect -270 -50 -225 -40
rect -205 -50 -195 20
rect -270 -60 -195 -50
rect -170 20 -130 30
rect -170 -50 -160 20
rect -140 -50 -130 20
rect -170 -60 -130 -50
rect -105 20 -65 30
rect -105 -50 -95 20
rect -75 -50 -65 20
rect 10 10 30 35
rect -105 -60 -65 -50
rect -15 0 135 10
rect -15 -10 105 0
rect -270 -255 -250 -60
rect -170 -85 -150 -60
rect -210 -105 -150 -85
rect -95 -85 -75 -60
rect -95 -105 -35 -85
rect -210 -125 -190 -105
rect -230 -135 -190 -125
rect -230 -205 -220 -135
rect -200 -205 -190 -135
rect -230 -215 -190 -205
rect -165 -135 -75 -125
rect -165 -205 -155 -135
rect -135 -205 -105 -135
rect -85 -205 -75 -135
rect -165 -215 -75 -205
rect -270 -265 -205 -255
rect -270 -275 -235 -265
rect -245 -335 -235 -275
rect -215 -335 -205 -265
rect -245 -345 -205 -335
rect -135 -265 -100 -255
rect -135 -335 -130 -265
rect -110 -325 -100 -265
rect -55 -265 -35 -105
rect -15 -90 5 -10
rect 95 -20 105 -10
rect 125 -20 135 0
rect 95 -30 135 -20
rect 30 -40 70 -30
rect 30 -60 40 -40
rect 60 -50 70 -40
rect 155 -50 175 35
rect 60 -60 175 -50
rect 30 -70 175 -60
rect 155 -90 175 -70
rect -15 -100 45 -90
rect -15 -110 15 -100
rect 5 -170 15 -110
rect 35 -170 45 -100
rect 5 -180 45 -170
rect 70 -100 110 -90
rect 70 -170 80 -100
rect 100 -170 110 -100
rect 70 -180 110 -170
rect 135 -100 175 -90
rect 135 -170 145 -100
rect 165 -170 175 -100
rect 135 -180 175 -170
rect 5 -200 25 -180
rect -15 -210 25 -200
rect -15 -230 -5 -210
rect 15 -230 25 -210
rect -15 -240 25 -230
rect 145 -255 165 -180
rect 35 -265 75 -255
rect -55 -285 45 -265
rect -25 -315 15 -305
rect -25 -325 -15 -315
rect -110 -335 -15 -325
rect 5 -335 15 -315
rect -135 -345 15 -335
rect 35 -335 45 -285
rect 65 -335 75 -265
rect 35 -345 75 -335
rect 145 -265 185 -255
rect 145 -335 155 -265
rect 175 -335 185 -265
rect 145 -345 185 -335
rect -180 -400 -140 -390
rect -180 -420 -170 -400
rect -150 -420 -140 -400
rect -180 -430 -140 -420
rect -80 -400 -40 -390
rect -80 -420 -70 -400
rect -50 -420 -40 -400
rect -80 -430 -40 -420
rect 75 -400 115 -390
rect 75 -420 85 -400
rect 105 -420 115 -400
rect 75 -430 115 -420
<< viali >>
rect -165 160 -145 230
rect 60 205 80 275
rect 110 205 130 275
rect -155 -205 -135 -135
rect -105 -205 -85 -135
rect 80 -170 100 -100
rect -170 -420 -150 -400
rect -70 -420 -50 -400
rect 85 -420 105 -400
<< metal1 >>
rect -275 275 205 415
rect -275 230 60 275
rect -275 160 -165 230
rect -145 205 60 230
rect 80 205 110 275
rect 130 205 205 275
rect -145 160 205 205
rect -275 150 205 160
rect 10 30 30 45
rect 155 30 175 35
rect -275 -100 205 30
rect -275 -135 80 -100
rect -275 -205 -155 -135
rect -135 -205 -105 -135
rect -85 -170 80 -135
rect 100 -170 205 -100
rect -85 -205 205 -170
rect -275 -345 205 -205
rect -275 -400 205 -390
rect -275 -420 -170 -400
rect -150 -420 -70 -400
rect -50 -420 85 -400
rect 105 -420 205 -400
rect -275 -430 205 -420
<< labels >>
rlabel metal1 -275 -410 -275 -410 7 clk
port 5 w
rlabel metal1 -275 -160 -275 -160 7 VN
port 4 w
rlabel locali -275 455 -275 455 7 D
port 1 w
rlabel metal1 -275 280 -275 280 7 VP
port 3 w
rlabel locali -275 400 -275 400 7 Dn
port 2 w
rlabel locali 205 400 205 400 3 Qn
port 7 e
rlabel locali 205 455 205 455 3 Q
port 6 e
<< end >>
