magic
tech sky130A
timestamp 1620681883
<< nwell >>
rect -100 435 300 535
<< nmos >>
rect -30 185 -15 360
rect 35 185 50 360
rect 100 185 115 360
rect 165 185 180 360
rect -85 90 265 105
<< pmos >>
rect -30 455 -15 515
rect 35 455 50 515
rect 100 455 115 515
rect 165 455 180 515
<< ndiff >>
rect -80 345 -30 360
rect -80 200 -65 345
rect -45 200 -30 345
rect -80 185 -30 200
rect -15 345 35 360
rect -15 200 0 345
rect 20 200 35 345
rect -15 185 35 200
rect 50 345 100 360
rect 50 200 65 345
rect 85 200 100 345
rect 50 185 100 200
rect 115 345 165 360
rect 115 200 130 345
rect 150 200 165 345
rect 115 185 165 200
rect 180 345 230 360
rect 180 200 195 345
rect 215 200 230 345
rect 180 185 230 200
rect -85 140 265 155
rect -85 120 -70 140
rect 250 120 265 140
rect -85 105 265 120
rect -85 75 265 90
rect -85 55 -70 75
rect 250 55 265 75
rect -85 40 265 55
<< pdiff >>
rect -80 500 -30 515
rect -80 470 -65 500
rect -45 470 -30 500
rect -80 455 -30 470
rect -15 500 35 515
rect -15 470 0 500
rect 20 470 35 500
rect -15 455 35 470
rect 50 500 100 515
rect 50 470 65 500
rect 85 470 100 500
rect 50 455 100 470
rect 115 500 165 515
rect 115 470 130 500
rect 150 470 165 500
rect 115 455 165 470
rect 180 500 230 515
rect 180 470 195 500
rect 215 470 230 500
rect 180 455 230 470
<< ndiffc >>
rect -65 200 -45 345
rect 0 200 20 345
rect 65 200 85 345
rect 130 200 150 345
rect 195 200 215 345
rect -70 120 250 140
rect -70 55 250 75
<< pdiffc >>
rect -65 470 -45 500
rect 0 470 20 500
rect 65 470 85 500
rect 130 470 150 500
rect 195 470 215 500
<< psubdiff >>
rect -85 25 265 40
rect -85 5 -70 25
rect 250 5 265 25
rect -85 -10 265 5
<< nsubdiff >>
rect 230 500 280 515
rect 230 470 245 500
rect 265 470 280 500
rect 230 455 280 470
<< psubdiffcont >>
rect -70 5 250 25
<< nsubdiffcont >>
rect 245 470 265 500
<< poly >>
rect -75 560 -35 570
rect -75 540 -65 560
rect -45 545 -35 560
rect 35 560 75 570
rect -45 540 -15 545
rect -75 530 -15 540
rect -30 515 -15 530
rect 35 540 45 560
rect 65 540 75 560
rect 185 560 225 570
rect 185 545 195 560
rect 35 530 75 540
rect 165 540 195 545
rect 215 540 225 560
rect 165 530 225 540
rect 35 515 50 530
rect 100 515 115 530
rect 165 515 180 530
rect -30 440 -15 455
rect -75 405 -35 415
rect -75 385 -65 405
rect -45 390 -35 405
rect -45 385 -15 390
rect -75 375 -15 385
rect -30 360 -15 375
rect 35 360 50 455
rect 100 435 115 455
rect 165 440 180 455
rect 75 425 115 435
rect 75 405 85 425
rect 105 405 115 425
rect 75 395 115 405
rect 100 360 115 395
rect 185 405 225 415
rect 185 390 195 405
rect 165 385 195 390
rect 215 385 225 405
rect 165 375 225 385
rect 165 360 180 375
rect -30 170 -15 185
rect 35 170 50 185
rect 100 170 115 185
rect 165 170 180 185
rect -100 90 -85 105
rect 265 90 300 105
<< polycont >>
rect -65 540 -45 560
rect 45 540 65 560
rect 195 540 215 560
rect -65 385 -45 405
rect 85 405 105 425
rect 195 385 215 405
<< locali >>
rect -75 560 -35 570
rect -75 540 -65 560
rect -45 540 -35 560
rect -75 530 -35 540
rect -65 510 -45 530
rect -10 510 10 590
rect 140 570 160 590
rect 35 560 160 570
rect 35 540 45 560
rect 65 550 160 560
rect 65 540 75 550
rect 35 530 75 540
rect 140 510 160 550
rect 185 560 225 570
rect 185 540 195 560
rect 215 540 225 560
rect 185 530 225 540
rect 195 510 215 530
rect -75 500 -35 510
rect -75 470 -65 500
rect -45 470 -35 500
rect -75 460 -35 470
rect -10 500 30 510
rect -10 470 0 500
rect 20 470 30 500
rect -10 460 30 470
rect 55 500 95 510
rect 55 470 65 500
rect 85 470 95 500
rect 55 460 95 470
rect 120 500 160 510
rect 120 470 130 500
rect 150 470 160 500
rect 120 460 160 470
rect 185 500 275 510
rect 185 470 195 500
rect 215 470 245 500
rect 265 470 275 500
rect 185 460 275 470
rect -10 415 10 460
rect 75 425 115 435
rect 75 415 85 425
rect -75 405 -35 415
rect -75 385 -65 405
rect -45 385 -35 405
rect -75 375 -35 385
rect -10 405 85 415
rect 105 405 115 425
rect -10 395 115 405
rect -65 355 -45 375
rect -10 355 10 395
rect 140 355 160 460
rect 185 405 225 415
rect 185 385 195 405
rect 215 385 225 405
rect 185 375 225 385
rect 195 355 215 375
rect -75 345 -35 355
rect -75 200 -65 345
rect -45 200 -35 345
rect -75 190 -35 200
rect -10 345 30 355
rect -10 200 0 345
rect 20 200 30 345
rect -10 190 30 200
rect 55 345 95 355
rect 55 200 65 345
rect 85 200 95 345
rect 55 150 95 200
rect 120 345 160 355
rect 120 200 130 345
rect 150 200 160 345
rect 120 190 160 200
rect 185 345 225 355
rect 185 200 195 345
rect 215 200 225 345
rect 185 190 225 200
rect -80 140 260 150
rect -80 120 -70 140
rect 250 120 260 140
rect -80 110 260 120
rect -80 75 260 85
rect -80 55 -70 75
rect 250 55 260 75
rect -80 25 260 55
rect -80 5 -70 25
rect 250 5 260 25
rect -80 -5 260 5
<< viali >>
rect -65 470 -45 500
rect 65 470 85 500
rect 195 470 215 500
rect 245 470 265 500
rect -70 55 250 75
rect -70 5 250 25
<< metal1 >>
rect -100 500 300 510
rect -100 470 -65 500
rect -45 470 65 500
rect 85 470 195 500
rect 215 470 245 500
rect 265 470 300 500
rect -100 460 300 470
rect -100 75 300 355
rect -100 55 -70 75
rect 250 55 300 75
rect -100 25 300 55
rect -100 5 -70 25
rect 250 5 300 25
rect -100 -5 300 5
<< labels >>
rlabel locali 150 590 150 590 1 Odd
rlabel locali 0 590 0 590 1 Even
rlabel metal1 -100 485 -100 485 7 VP
rlabel metal1 -100 185 -100 185 7 VN
rlabel poly -100 95 -100 95 7 En
<< end >>
