magic
tech sky130A
timestamp 1620496349
<< error_p >>
rect -71 338 -65 341
rect -21 338 -15 341
rect 214 338 220 341
rect 314 338 320 341
rect -88 335 -62 338
rect -38 335 -12 338
rect 197 335 223 338
rect 297 335 323 338
rect -91 332 -59 335
rect -91 329 -82 332
rect -85 18 -82 329
rect -68 329 -59 332
rect -41 332 -9 335
rect -41 329 -32 332
rect -68 18 -62 329
rect -85 15 -62 18
rect -35 18 -32 329
rect -18 329 -9 332
rect 194 332 226 335
rect 194 329 203 332
rect -18 18 -12 329
rect 200 308 203 329
rect 217 329 226 332
rect 294 332 326 335
rect 294 329 303 332
rect 217 308 223 329
rect 200 305 223 308
rect 300 308 303 329
rect 317 329 326 332
rect 317 308 323 329
rect 300 305 323 308
rect 214 302 223 305
rect 314 302 323 305
rect 214 299 220 302
rect 314 299 320 302
rect -35 15 -12 18
rect -71 12 -62 15
rect -21 12 -12 15
rect -71 9 -65 12
rect -21 9 -15 12
<< nwell >>
rect 100 270 420 370
<< nmos >>
rect 0 0 15 350
rect 170 40 185 215
rect 235 40 250 215
<< pmos >>
rect 170 290 185 350
rect 335 290 350 350
<< ndiff >>
rect -50 335 0 350
rect -50 15 -35 335
rect -15 15 0 335
rect -50 0 0 15
rect 15 335 65 350
rect 15 15 30 335
rect 50 15 65 335
rect 120 200 170 215
rect 120 55 135 200
rect 155 55 170 200
rect 120 40 170 55
rect 185 200 235 215
rect 185 55 200 200
rect 220 55 235 200
rect 185 40 235 55
rect 250 200 300 215
rect 250 55 265 200
rect 285 55 300 200
rect 250 40 300 55
rect 15 0 65 15
<< pdiff >>
rect 120 335 170 350
rect 120 305 135 335
rect 155 305 170 335
rect 120 290 170 305
rect 185 335 235 350
rect 285 335 335 350
rect 185 305 200 335
rect 220 305 235 335
rect 285 305 300 335
rect 320 305 335 335
rect 185 290 235 305
rect 285 290 335 305
rect 350 335 400 350
rect 350 305 365 335
rect 385 305 400 335
rect 350 290 400 305
<< ndiffc >>
rect -35 15 -15 335
rect 30 15 50 335
rect 135 55 155 200
rect 200 55 220 200
rect 265 55 285 200
<< pdiffc >>
rect 135 305 155 335
rect 200 305 220 335
rect 300 305 320 335
rect 365 305 385 335
<< psubdiff >>
rect -100 335 -50 350
rect -100 15 -85 335
rect -65 15 -50 335
rect -100 0 -50 15
<< nsubdiff >>
rect 235 335 285 350
rect 235 305 250 335
rect 270 305 285 335
rect 235 290 285 305
<< psubdiffcont >>
rect -85 15 -65 335
<< nsubdiffcont >>
rect 250 305 270 335
<< poly >>
rect 310 435 350 445
rect 310 415 320 435
rect 340 415 350 435
rect 310 405 350 415
rect 170 395 210 405
rect 170 375 180 395
rect 200 375 210 395
rect 170 365 210 375
rect 0 350 15 365
rect 170 350 185 365
rect 335 350 350 405
rect 170 215 185 290
rect 215 265 255 270
rect 335 265 350 290
rect 215 260 350 265
rect 215 240 225 260
rect 245 250 350 260
rect 245 240 255 250
rect 215 230 255 240
rect 235 215 250 230
rect 170 25 185 40
rect 235 25 250 40
rect 0 -15 15 0
<< polycont >>
rect 320 415 340 435
rect 180 375 200 395
rect 225 240 245 260
<< locali >>
rect 170 405 190 465
rect 330 445 350 465
rect 310 435 350 445
rect 310 415 320 435
rect 340 415 350 435
rect 310 405 350 415
rect 170 395 210 405
rect 170 375 180 395
rect 200 385 210 395
rect 200 375 375 385
rect 170 365 375 375
rect 355 345 375 365
rect -95 335 -5 345
rect -95 15 -85 335
rect -65 15 -35 335
rect -15 15 -5 335
rect -95 5 -5 15
rect 20 335 60 345
rect 20 15 30 335
rect 50 25 60 335
rect 125 335 165 345
rect 125 305 135 335
rect 155 305 165 335
rect 125 295 165 305
rect 190 335 330 345
rect 190 305 200 335
rect 220 305 250 335
rect 270 305 300 335
rect 320 305 330 335
rect 190 295 330 305
rect 355 335 395 345
rect 355 305 365 335
rect 385 305 395 335
rect 355 295 395 305
rect 135 270 155 295
rect 135 260 255 270
rect 135 250 225 260
rect 135 210 155 250
rect 215 240 225 250
rect 245 240 255 260
rect 215 230 255 240
rect 355 210 375 295
rect 125 200 165 210
rect 125 55 135 200
rect 155 55 165 200
rect 125 45 165 55
rect 190 200 230 210
rect 190 55 200 200
rect 220 55 230 200
rect 190 45 230 55
rect 255 200 375 210
rect 255 55 265 200
rect 285 190 375 200
rect 285 55 295 190
rect 255 45 295 55
rect 190 25 210 45
rect 50 15 210 25
rect 20 5 210 15
<< viali >>
rect -85 15 -65 335
rect -35 15 -15 335
rect 200 305 220 335
rect 300 305 320 335
<< end >>
