magic
tech sky130A
timestamp 1620748619
<< nwell >>
rect -430 480 280 920
<< nmos >>
rect -360 200 -345 400
rect -295 200 -280 400
rect -230 200 -215 400
rect -165 200 -150 400
rect 0 200 15 400
rect 65 200 80 400
rect 130 200 145 400
rect 195 200 210 400
<< pmos >>
rect -360 500 -345 900
rect -295 500 -280 900
rect -230 500 -215 900
rect -165 500 -150 900
rect 0 500 15 900
rect 65 500 80 900
rect 130 500 145 900
rect 195 500 210 900
<< ndiff >>
rect -410 385 -360 400
rect -410 215 -395 385
rect -375 215 -360 385
rect -410 200 -360 215
rect -345 385 -295 400
rect -345 215 -330 385
rect -310 215 -295 385
rect -345 200 -295 215
rect -280 385 -230 400
rect -280 215 -265 385
rect -245 215 -230 385
rect -280 200 -230 215
rect -215 385 -165 400
rect -215 215 -200 385
rect -180 215 -165 385
rect -215 200 -165 215
rect -150 385 -100 400
rect -50 385 0 400
rect -150 215 -135 385
rect -115 215 -100 385
rect -50 215 -35 385
rect -15 215 0 385
rect -150 200 -100 215
rect -50 200 0 215
rect 15 385 65 400
rect 15 215 30 385
rect 50 215 65 385
rect 15 200 65 215
rect 80 385 130 400
rect 80 215 95 385
rect 115 215 130 385
rect 80 200 130 215
rect 145 385 195 400
rect 145 215 160 385
rect 180 215 195 385
rect 145 200 195 215
rect 210 385 260 400
rect 210 215 225 385
rect 245 215 260 385
rect 210 200 260 215
<< pdiff >>
rect -410 885 -360 900
rect -410 515 -395 885
rect -375 515 -360 885
rect -410 500 -360 515
rect -345 885 -295 900
rect -345 515 -330 885
rect -310 515 -295 885
rect -345 500 -295 515
rect -280 885 -230 900
rect -280 515 -265 885
rect -245 515 -230 885
rect -280 500 -230 515
rect -215 885 -165 900
rect -215 515 -200 885
rect -180 515 -165 885
rect -215 500 -165 515
rect -150 885 -100 900
rect -50 885 0 900
rect -150 515 -135 885
rect -115 515 -100 885
rect -50 515 -35 885
rect -15 515 0 885
rect -150 500 -100 515
rect -50 500 0 515
rect 15 885 65 900
rect 15 515 30 885
rect 50 515 65 885
rect 15 500 65 515
rect 80 885 130 900
rect 80 515 95 885
rect 115 515 130 885
rect 80 500 130 515
rect 145 885 195 900
rect 145 515 160 885
rect 180 515 195 885
rect 145 500 195 515
rect 210 885 260 900
rect 210 515 225 885
rect 245 515 260 885
rect 210 500 260 515
<< ndiffc >>
rect -395 215 -375 385
rect -330 215 -310 385
rect -265 215 -245 385
rect -200 215 -180 385
rect -135 215 -115 385
rect -35 215 -15 385
rect 30 215 50 385
rect 95 215 115 385
rect 160 215 180 385
rect 225 215 245 385
<< pdiffc >>
rect -395 515 -375 885
rect -330 515 -310 885
rect -265 515 -245 885
rect -200 515 -180 885
rect -135 515 -115 885
rect -35 515 -15 885
rect 30 515 50 885
rect 95 515 115 885
rect 160 515 180 885
rect 225 515 245 885
<< psubdiff >>
rect -100 385 -50 400
rect -100 215 -85 385
rect -65 215 -50 385
rect -100 200 -50 215
<< nsubdiff >>
rect -100 885 -50 900
rect -100 515 -85 885
rect -65 515 -50 885
rect -100 500 -50 515
<< psubdiffcont >>
rect -85 215 -65 385
<< nsubdiffcont >>
rect -85 515 -65 885
<< poly >>
rect -400 945 -360 955
rect -400 925 -390 945
rect -370 930 -360 945
rect -95 945 -55 955
rect -95 930 -85 945
rect -370 925 -345 930
rect -400 915 -345 925
rect -165 925 -85 930
rect -65 930 -55 945
rect -65 925 15 930
rect -165 915 15 925
rect -360 900 -345 915
rect -295 900 -280 915
rect -230 900 -215 915
rect -165 900 -150 915
rect 0 900 15 915
rect 65 900 80 915
rect 130 900 145 915
rect 195 900 210 915
rect -360 485 -345 500
rect -400 445 -360 455
rect -400 425 -390 445
rect -370 430 -360 445
rect -370 425 -345 430
rect -400 415 -345 425
rect -360 400 -345 415
rect -295 400 -280 500
rect -230 400 -215 500
rect -165 485 -150 500
rect 0 485 15 500
rect -95 445 -55 455
rect -95 430 -85 445
rect -165 425 -85 430
rect -65 430 -55 445
rect -65 425 15 430
rect -165 415 15 425
rect -165 400 -150 415
rect 0 400 15 415
rect 65 400 80 500
rect 130 400 145 500
rect 195 485 210 500
rect 195 475 250 485
rect 195 470 220 475
rect 210 455 220 470
rect 240 455 250 475
rect 210 445 250 455
rect 195 400 210 415
rect -360 185 -345 200
rect -295 185 -280 200
rect -230 185 -215 200
rect -165 185 -150 200
rect 0 185 15 200
rect 65 185 80 200
rect 130 185 145 200
rect 195 185 210 200
rect -295 175 -255 185
rect -295 155 -285 175
rect -265 155 -255 175
rect -295 145 -255 155
rect -230 175 -190 185
rect -230 155 -220 175
rect -200 155 -190 175
rect -230 145 -190 155
rect 65 175 105 185
rect 65 155 75 175
rect 95 155 105 175
rect 65 145 105 155
rect 130 175 170 185
rect 130 155 140 175
rect 160 155 170 175
rect 195 175 250 185
rect 195 170 220 175
rect 130 145 170 155
rect 210 155 220 170
rect 240 155 250 175
rect 210 145 250 155
<< polycont >>
rect -390 925 -370 945
rect -85 925 -65 945
rect -390 425 -370 445
rect -85 425 -65 445
rect 220 455 240 475
rect -285 155 -265 175
rect -220 155 -200 175
rect 75 155 95 175
rect 140 155 160 175
rect 220 155 240 175
<< locali >>
rect -330 1040 280 1060
rect -400 945 -360 955
rect -400 925 -390 945
rect -370 925 -360 945
rect -400 915 -360 925
rect -395 895 -375 915
rect -330 895 -310 1040
rect -200 1000 280 1020
rect -200 895 -180 1000
rect 30 960 280 980
rect -95 945 -55 955
rect -95 925 -85 945
rect -65 925 -55 945
rect -95 895 -55 925
rect 30 895 50 960
rect 160 920 280 940
rect 160 895 180 920
rect -405 885 -360 895
rect -405 515 -395 885
rect -375 515 -360 885
rect -405 505 -360 515
rect -340 885 -295 895
rect -340 515 -330 885
rect -310 515 -295 885
rect -340 505 -295 515
rect -275 885 -230 895
rect -275 515 -265 885
rect -245 515 -230 885
rect -275 505 -230 515
rect -210 885 -165 895
rect -210 515 -200 885
rect -180 515 -165 885
rect -210 505 -165 515
rect -145 885 -5 895
rect -145 515 -135 885
rect -115 515 -85 885
rect -65 515 -35 885
rect -15 515 -5 885
rect -145 505 -5 515
rect 20 885 60 895
rect 20 515 30 885
rect 50 515 60 885
rect 20 505 60 515
rect 85 885 125 895
rect 85 515 95 885
rect 115 515 125 885
rect 85 505 125 515
rect 150 885 190 895
rect 150 515 160 885
rect 180 515 190 885
rect 150 505 190 515
rect 215 885 255 895
rect 215 515 225 885
rect 245 515 255 885
rect 215 505 255 515
rect -400 445 -360 455
rect -400 425 -390 445
rect -370 425 -360 445
rect -400 415 -360 425
rect -395 395 -375 415
rect -330 395 -310 505
rect -200 395 -180 505
rect -95 445 -55 455
rect -95 425 -85 445
rect -65 425 -55 445
rect -95 395 -55 425
rect 30 395 50 505
rect 160 395 180 505
rect 225 485 245 505
rect 210 475 250 485
rect 210 455 220 475
rect 240 455 250 475
rect 210 445 250 455
rect -405 385 -360 395
rect -405 215 -395 385
rect -375 215 -360 385
rect -405 205 -360 215
rect -340 385 -295 395
rect -340 215 -330 385
rect -310 215 -295 385
rect -340 205 -295 215
rect -275 385 -230 395
rect -275 215 -265 385
rect -245 215 -230 385
rect -275 205 -230 215
rect -210 385 -165 395
rect -210 215 -200 385
rect -180 215 -165 385
rect -210 205 -165 215
rect -145 385 -5 395
rect -145 215 -135 385
rect -115 215 -85 385
rect -65 215 -35 385
rect -15 215 -5 385
rect -145 205 -5 215
rect 20 385 60 395
rect 20 215 30 385
rect 50 215 60 385
rect 20 205 60 215
rect 85 385 125 395
rect 85 215 95 385
rect 115 215 125 385
rect 85 205 125 215
rect 150 385 190 395
rect 150 215 160 385
rect 180 215 190 385
rect 150 205 190 215
rect 215 385 255 395
rect 215 215 225 385
rect 245 215 255 385
rect 215 205 255 215
rect 225 185 245 205
rect -295 175 -255 185
rect -295 165 -285 175
rect -430 155 -285 165
rect -265 155 -255 175
rect -430 145 -255 155
rect -230 175 -190 185
rect -230 155 -220 175
rect -200 155 -190 175
rect -230 145 -190 155
rect 65 175 105 185
rect 65 155 75 175
rect 95 155 105 175
rect 65 145 105 155
rect 130 175 170 185
rect 130 155 140 175
rect 160 155 170 175
rect 130 145 170 155
rect 210 175 250 185
rect 210 155 220 175
rect 240 155 250 175
rect 210 145 250 155
rect -230 125 -210 145
rect -430 105 -210 125
rect 65 85 85 145
rect -430 65 85 85
rect 130 45 150 145
rect -430 25 150 45
<< viali >>
rect -395 515 -375 885
rect -265 515 -245 885
rect -135 515 -115 885
rect -85 515 -65 885
rect -35 515 -15 885
rect 95 515 115 885
rect 225 515 245 885
rect -395 215 -375 385
rect -265 215 -245 385
rect -135 215 -115 385
rect -85 215 -65 385
rect -35 215 -15 385
rect 95 215 115 385
rect 225 215 245 385
<< metal1 >>
rect -430 885 280 895
rect -430 515 -395 885
rect -375 515 -265 885
rect -245 515 -135 885
rect -115 515 -85 885
rect -65 515 -35 885
rect -15 515 95 885
rect 115 515 225 885
rect 245 515 280 885
rect -430 505 280 515
rect -430 385 280 395
rect -430 215 -395 385
rect -375 215 -265 385
rect -245 215 -135 385
rect -115 215 -85 385
rect -65 215 -35 385
rect -15 215 95 385
rect 115 215 225 385
rect 245 215 280 385
rect -430 205 280 215
<< labels >>
rlabel locali 280 1050 280 1050 3 Q0
rlabel locali 280 1010 280 1010 3 Q1
rlabel locali 280 970 280 970 3 Q2
rlabel locali 280 930 280 930 3 Q3
rlabel metal1 -430 685 -430 685 7 VP
rlabel metal1 -430 310 -430 310 7 VN
rlabel locali -430 155 -430 155 7 A0A1
rlabel locali -430 115 -430 115 7 A0nA1
rlabel locali -430 75 -430 75 7 A0A1n
rlabel locali -430 35 -430 35 7 A0nA1n
<< end >>
