magic
tech sky130A
timestamp 1620758043
<< error_p >>
rect -526 88 -520 91
rect -476 88 -470 91
rect -411 88 -405 91
rect -281 88 -275 91
rect -151 88 -145 91
rect -21 88 -15 91
rect 109 88 115 91
rect 174 88 180 91
rect -543 85 -517 88
rect -493 85 -467 88
rect -428 85 -402 88
rect -298 85 -272 88
rect -168 85 -142 88
rect -38 85 -12 88
rect 92 85 118 88
rect 157 85 183 88
rect -546 82 -514 85
rect -546 79 -537 82
rect -540 18 -537 79
rect -523 79 -514 82
rect -496 82 -464 85
rect -496 79 -487 82
rect -523 18 -517 79
rect -540 15 -517 18
rect -490 18 -487 79
rect -473 79 -464 82
rect -431 82 -399 85
rect -431 79 -422 82
rect -473 18 -467 79
rect -490 15 -467 18
rect -425 18 -422 79
rect -408 79 -399 82
rect -301 82 -269 85
rect -301 79 -292 82
rect -408 18 -402 79
rect -425 15 -402 18
rect -295 18 -292 79
rect -278 79 -269 82
rect -171 82 -139 85
rect -171 79 -162 82
rect -278 18 -272 79
rect -295 15 -272 18
rect -165 18 -162 79
rect -148 79 -139 82
rect -41 82 -9 85
rect -41 79 -32 82
rect -148 18 -142 79
rect -165 15 -142 18
rect -35 18 -32 79
rect -18 79 -9 82
rect 89 82 121 85
rect 89 79 98 82
rect -18 18 -12 79
rect -35 15 -12 18
rect 95 18 98 79
rect 112 79 121 82
rect 154 82 186 85
rect 154 79 163 82
rect 112 18 118 79
rect 95 15 118 18
rect 160 18 163 79
rect 177 79 186 82
rect 177 18 183 79
rect 160 15 183 18
rect -526 12 -517 15
rect -476 12 -467 15
rect -411 12 -402 15
rect -281 12 -272 15
rect -151 12 -142 15
rect -21 12 -12 15
rect 109 12 118 15
rect 174 12 183 15
rect -526 9 -520 12
rect -476 9 -470 12
rect -411 9 -405 12
rect -281 9 -275 12
rect -151 9 -145 12
rect -21 9 -15 12
rect 109 9 115 12
rect 174 9 180 12
<< nmos >>
rect -455 200 -440 400
rect -390 200 -375 400
rect -325 200 -310 400
rect -260 200 -245 400
rect 45 200 60 400
rect 110 200 125 400
rect 175 200 190 400
rect 240 200 255 400
rect -455 0 -440 100
rect -390 0 -375 100
rect -325 0 -310 100
rect -260 0 -245 100
rect -195 0 -180 100
rect -130 0 -115 100
rect -65 0 -50 100
rect 0 0 15 100
rect 65 0 80 100
rect 130 0 145 100
<< ndiff >>
rect -505 385 -455 400
rect -505 215 -490 385
rect -470 215 -455 385
rect -505 200 -455 215
rect -440 385 -390 400
rect -440 215 -425 385
rect -405 215 -390 385
rect -440 200 -390 215
rect -375 385 -325 400
rect -375 215 -360 385
rect -340 215 -325 385
rect -375 200 -325 215
rect -310 385 -260 400
rect -310 215 -295 385
rect -275 215 -260 385
rect -310 200 -260 215
rect -245 385 -195 400
rect -245 215 -230 385
rect -210 215 -195 385
rect -245 200 -195 215
rect -5 385 45 400
rect -5 215 10 385
rect 30 215 45 385
rect -5 200 45 215
rect 60 385 110 400
rect 60 215 75 385
rect 95 215 110 385
rect 60 200 110 215
rect 125 385 175 400
rect 125 215 140 385
rect 160 215 175 385
rect 125 200 175 215
rect 190 385 240 400
rect 190 215 205 385
rect 225 215 240 385
rect 190 200 240 215
rect 255 385 305 400
rect 255 215 270 385
rect 290 215 305 385
rect 255 200 305 215
rect -505 85 -455 100
rect -505 15 -490 85
rect -470 15 -455 85
rect -505 0 -455 15
rect -440 85 -390 100
rect -440 15 -425 85
rect -405 15 -390 85
rect -440 0 -390 15
rect -375 85 -325 100
rect -375 15 -360 85
rect -340 15 -325 85
rect -375 0 -325 15
rect -310 85 -260 100
rect -310 15 -295 85
rect -275 15 -260 85
rect -310 0 -260 15
rect -245 85 -195 100
rect -245 15 -230 85
rect -210 15 -195 85
rect -245 0 -195 15
rect -180 85 -130 100
rect -180 15 -165 85
rect -145 15 -130 85
rect -180 0 -130 15
rect -115 85 -65 100
rect -115 15 -100 85
rect -80 15 -65 85
rect -115 0 -65 15
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 145 85 195 100
rect 145 15 160 85
rect 180 15 195 85
rect 145 0 195 15
<< ndiffc >>
rect -490 215 -470 385
rect -425 215 -405 385
rect -360 215 -340 385
rect -295 215 -275 385
rect -230 215 -210 385
rect 10 215 30 385
rect 75 215 95 385
rect 140 215 160 385
rect 205 215 225 385
rect 270 215 290 385
rect -490 15 -470 85
rect -425 15 -405 85
rect -360 15 -340 85
rect -295 15 -275 85
rect -230 15 -210 85
rect -165 15 -145 85
rect -100 15 -80 85
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
rect 160 15 180 85
<< psubdiff >>
rect -555 385 -505 400
rect -555 215 -540 385
rect -520 215 -505 385
rect -555 200 -505 215
rect -55 385 -5 400
rect -55 215 -40 385
rect -20 215 -5 385
rect -55 200 -5 215
rect -555 85 -505 100
rect -555 15 -540 85
rect -520 15 -505 85
rect -555 0 -505 15
<< psubdiffcont >>
rect -540 215 -520 385
rect -40 215 -20 385
rect -540 15 -520 85
<< poly >>
rect -455 400 -440 415
rect -390 400 -375 415
rect -325 400 -310 415
rect -260 400 -245 415
rect 45 400 60 415
rect 110 400 125 415
rect 175 400 190 415
rect 240 400 255 415
rect -455 185 -440 200
rect -390 185 -375 200
rect -325 185 -310 200
rect -260 185 -245 200
rect 45 185 60 200
rect 110 185 125 200
rect 175 185 190 200
rect 240 185 255 200
rect -495 145 -455 155
rect -495 125 -485 145
rect -465 130 -455 145
rect -465 125 -440 130
rect -495 115 -440 125
rect -455 100 -440 115
rect -390 100 -375 115
rect -325 100 -310 115
rect -260 100 -245 115
rect -195 100 -180 115
rect -130 100 -115 115
rect -65 100 -50 115
rect 0 100 15 115
rect 65 100 80 115
rect 130 100 145 115
rect -455 -15 -440 0
rect -390 -15 -375 0
rect -325 -15 -310 0
rect -260 -15 -245 0
rect -195 -15 -180 0
rect -130 -15 -115 0
rect -65 -15 -50 0
rect 0 -15 15 0
rect 65 -15 80 0
rect 130 -15 145 0
rect 130 -25 185 -15
rect 130 -30 155 -25
rect 145 -45 155 -30
rect 175 -45 185 -25
rect 145 -55 185 -45
<< polycont >>
rect -485 125 -465 145
rect 155 -45 175 -25
<< locali >>
rect -550 385 -460 395
rect -550 215 -540 385
rect -520 215 -490 385
rect -470 215 -460 385
rect -550 205 -460 215
rect -440 385 -395 395
rect -440 215 -425 385
rect -405 215 -395 385
rect -440 205 -395 215
rect -375 385 -330 395
rect -375 215 -360 385
rect -340 215 -330 385
rect -375 205 -330 215
rect -310 385 -265 395
rect -310 215 -295 385
rect -275 215 -265 385
rect -310 205 -265 215
rect -245 385 -200 395
rect -245 215 -230 385
rect -210 215 -200 385
rect -245 205 -200 215
rect -50 385 40 395
rect -50 215 -40 385
rect -20 215 10 385
rect 30 215 40 385
rect -50 205 40 215
rect 60 385 105 395
rect 60 215 75 385
rect 95 215 105 385
rect 60 205 105 215
rect 125 385 170 395
rect 125 215 140 385
rect 160 215 170 385
rect 125 205 170 215
rect 190 385 235 395
rect 190 215 205 385
rect 225 215 235 385
rect 190 205 235 215
rect 255 385 300 395
rect 255 215 270 385
rect 290 215 300 385
rect 255 205 300 215
rect -495 145 -455 155
rect -495 125 -485 145
rect -465 125 -455 145
rect -495 115 -455 125
rect -490 95 -470 115
rect -550 85 -460 95
rect -550 15 -540 85
rect -520 15 -490 85
rect -470 15 -460 85
rect -550 5 -460 15
rect -435 85 -395 95
rect -435 15 -425 85
rect -405 15 -395 85
rect -435 5 -395 15
rect -370 85 -330 95
rect -370 15 -360 85
rect -340 15 -330 85
rect -370 5 -330 15
rect -305 85 -265 95
rect -305 15 -295 85
rect -275 15 -265 85
rect -305 5 -265 15
rect -240 85 -200 95
rect -240 15 -230 85
rect -210 15 -200 85
rect -240 5 -200 15
rect -175 85 -135 95
rect -175 15 -165 85
rect -145 15 -135 85
rect -175 5 -135 15
rect -110 85 -70 95
rect -110 15 -100 85
rect -80 15 -70 85
rect -110 5 -70 15
rect -45 85 -5 95
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 5 -5 15
rect 20 85 60 95
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect 85 5 125 15
rect 150 85 190 95
rect 150 15 160 85
rect 180 15 190 85
rect 150 5 190 15
rect 160 -15 180 5
rect 145 -25 185 -15
rect 145 -45 155 -25
rect 175 -45 185 -25
rect 145 -55 185 -45
<< viali >>
rect -540 15 -520 85
rect -490 15 -470 85
rect -425 15 -405 85
rect -295 15 -275 85
rect -165 15 -145 85
rect -35 15 -15 85
rect 95 15 115 85
rect 160 15 180 85
<< end >>
